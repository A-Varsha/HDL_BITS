module top_module (
    output out);
    wire  gnd;
assign out = gnd;
endmodule
